b0VIM 8.0      8�]t  v  leeunx                                  leeunx-VirtualBox                       ~leeunx/Algorithms/C/LongestIncreasingSubsequence/LongestIncreasingSubsequence.c                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           *                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             ad  Q       *       �  �  �  �  �  |  ^  F    �  �  �  �  c  a  `  >  )      �  �  �  �  l  :    �  �  �  �  �  �  |  q  d  b  a  U  4                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         } 	printf("%d", LIS(nums, 5)); 	int nums[5] = {0, 8, 4, 12, 3}; int main(){  } 	return len; 	puts(""); 		printf("%d ", dp[i]); 	for( int i = 0; i < length; i++ ) 	} 		printf("len: %d\n", len); 		if( index == len )len++;                  puts("");                         printf("%d ", dp[i]);                 for( int i = 0; i < length; i++ ) 		dp[index] = nums[num]; 	     	printf("%d\n", index); 		index = binarysearch(dp, 0, len, nums[num] ); 	for(int num = 0; num < length; num++){ 	dp = (int*)malloc(length);         	int* dp; 	int len = 0, index; int LIS( int* nums, int length ){  }         return (low + high)/2;  	printf("low: %d, high: %d\n", low, high);         }                 else low = mid + 1;                 else if( dp[mid] < num ) high = mid - 1;                 if( dp[mid] == num ) return mid; 		mid = (low + high)/2;         while( low <= high ){         int mid; int binarysearch(int* dp, int low, int high, int num){  #include <string.h> #include <stdlib.h> #include <stdio.h> 